// Copyright (C) 2023 Alan Jian (alanjian85@outlook.com)
// SPDX-License-Identifier: GPL-3.0

(* use_dsp = "yes" *) module rasterizer(
        input [9:0] x,
        input [9:0] y,
        output [19:0] ua,
        output [19:0] va,
        output [19:0] wa,
        output [19:0] a,
        output visible
    );

    localparam AX = 320;
    localparam AY = 60;

    localparam BX = 112;
    localparam BY = 420;
    localparam ABX = BX - AX;
    localparam ABY = BY - AY;

    localparam CX = 528;
    localparam CY = 420;
    localparam ACX = CX - AX;
    localparam ACY = CY - AY;

    localparam ABXACY = ABX * ACY;
    localparam ABYACX = ABY * ACX;
    localparam SA = ABXACY - ABYACX;
    assign a = SA > 0 ? SA : -SA;

    wire signed [9:0] apx = x - AX;
    wire signed [9:0] apy = y - AY;

    wire signed [19:0] abxapy = ABX * apy;
    wire signed [19:0] abyapx = ABY * apx;
    assign va = SA > 0 ? abxapy - abyapx : abyapx - abxapy;

    wire signed [19:0] apxacy = apx * ACY;
    wire signed [19:0] apyacx = apy * ACX;
    assign wa = SA > 0 ? apxacy - apyacx : apyacx - apxacy;

    assign ua = a - va - wa;

    assign visible = !(ua[19] || va[19] || wa[19]);

endmodule
