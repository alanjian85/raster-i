module top(
    input clk,
    input resetn,
    output [13:0] ddr3_addr,
    output [2:0]  ddr3_ba,
    output ddr3_cas_n,
    output [0:0]  ddr3_ck_n,
    output [0:0]  ddr3_ck_p,
    output [0:0]  ddr3_cke,
    output [0:0]  ddr3_cs_n,
    output [1:0]  ddr3_dm,
    inout  [15:0] ddr3_dq,
    inout  [1:0]  ddr3_dqs_n,
    inout  [1:0]  ddr3_dqs_p,
    output [0:0]  ddr3_odt,
    output ddr3_ras_n,
    output ddr3_reset_n,
    output ddr3_we_n,
    output [3:0] vga_r,
    output [3:0] vga_g,
    output [3:0] vga_b,
    output vga_hsync,
    output vga_vsync
);
    Trinity trinity(
        .clock(clk),
        .reset(!resetn),
        .io_ddr3_addr(ddr3_addr),
        .io_ddr3_ba(ddr3_ba),
        .io_ddr3_cas_n(ddr3_cas_n),
        .io_ddr3_ck_n(ddr3_ck_n),
        .io_ddr3_ck_p(ddr3_ck_p),
        .io_ddr3_cke(ddr3_cke),
        .io_ddr3_cs_n(ddr3_cs_n),
        .io_ddr3_dm(ddr3_dm),
        .io_ddr3_dq(ddr3_dq),
        .io_ddr3_dqs_n(ddr3_dqs_n),
        .io_ddr3_dqs_p(ddr3_dqs_p),
        .io_ddr3_odt(ddr3_odt),
        .io_ddr3_ras_n(ddr3_ras_n),
        .io_ddr3_reset_n(ddr3_reset_n),
        .io_ddr3_we_n(ddr3_we_n),
        .io_vga_r(vga_r),
        .io_vga_g(vga_g),
        .io_vga_b(vga_b),
        .io_vga_hsync(vga_hsync),
        .io_vga_vsync(vga_vsync)
    );
endmodule